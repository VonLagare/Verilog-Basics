module display ();

$display(& 1'b10);

$display(| 3'b101x);

$display(^ 4'b1101);


endmodule